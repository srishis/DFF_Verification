class dff_env;

	// instantiate all classes in environment
	dff_generator gen;
	dff_driver drv;
	dff_monitor mon;
	dff_coverage cov;
	dff_scoreboard sb;
	dff_ref_model rm;
	
	// create object for all classes
	function new();
		gen =	new();
		drv =	new();
		mon =	new();
		cov =	new();
		sb  =	new();
		rm  =   new();
	endfunction

	// call all run methods of each call in fork-join_none
	task run();
		fork
		gen.run();
		drv.run();
		mon.run();
		cov.run();
		sb.run();
		rm.run();
		join_none
	endtask

	task report();
		if(dff_cfg::error_count == 0)
			$display("Test failed with errors = %d", dff_cfg::error_count);
		else
			$display("TEST PASS: DFF Works as expected!!!");		
	endtask
	
endclass
