class dff_sb;
endclass