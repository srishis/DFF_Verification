class dff_golden;









endclass